module top (out,n9,n10,n13,n14,n16,n17,n24,n25,n27
        ,n28,n30,n36,n40,n43,n63,n173,n176,n178,n185
        ,n187,n194,n198,n219);
output out;
input n9;
input n10;
input n13;
input n14;
input n16;
input n17;
input n24;
input n25;
input n27;
input n28;
input n30;
input n36;
input n40;
input n43;
input n63;
input n173;
input n176;
input n178;
input n185;
input n187;
input n194;
input n198;
input n219;
wire n0;
wire n1;
wire n2;
wire n3;
wire n4;
wire n5;
wire n6;
wire n7;
wire n8;
wire n11;
wire n12;
wire n15;
wire n18;
wire n19;
wire n20;
wire n21;
wire n22;
wire n23;
wire n26;
wire n29;
wire n31;
wire n32;
wire n33;
wire n34;
wire n35;
wire n37;
wire n38;
wire n39;
wire n41;
wire n42;
wire n44;
wire n45;
wire n46;
wire n47;
wire n48;
wire n49;
wire n50;
wire n51;
wire n52;
wire n53;
wire n54;
wire n55;
wire n56;
wire n57;
wire n58;
wire n59;
wire n60;
wire n61;
wire n62;
wire n64;
wire n65;
wire n66;
wire n67;
wire n68;
wire n69;
wire n70;
wire n71;
wire n72;
wire n73;
wire n74;
wire n75;
wire n76;
wire n77;
wire n78;
wire n79;
wire n80;
wire n81;
wire n82;
wire n83;
wire n84;
wire n85;
wire n86;
wire n87;
wire n88;
wire n89;
wire n90;
wire n91;
wire n92;
wire n93;
wire n94;
wire n95;
wire n96;
wire n97;
wire n98;
wire n99;
wire n100;
wire n101;
wire n102;
wire n103;
wire n104;
wire n105;
wire n106;
wire n107;
wire n108;
wire n109;
wire n110;
wire n111;
wire n112;
wire n113;
wire n114;
wire n115;
wire n116;
wire n117;
wire n118;
wire n119;
wire n120;
wire n121;
wire n122;
wire n123;
wire n124;
wire n125;
wire n126;
wire n127;
wire n128;
wire n129;
wire n130;
wire n131;
wire n132;
wire n133;
wire n134;
wire n135;
wire n136;
wire n137;
wire n138;
wire n139;
wire n140;
wire n141;
wire n142;
wire n143;
wire n144;
wire n145;
wire n146;
wire n147;
wire n148;
wire n149;
wire n150;
wire n151;
wire n152;
wire n153;
wire n154;
wire n155;
wire n156;
wire n157;
wire n158;
wire n159;
wire n160;
wire n161;
wire n162;
wire n163;
wire n164;
wire n165;
wire n166;
wire n167;
wire n168;
wire n169;
wire n170;
wire n171;
wire n172;
wire n174;
wire n175;
wire n177;
wire n179;
wire n180;
wire n181;
wire n182;
wire n183;
wire n184;
wire n186;
wire n188;
wire n189;
wire n190;
wire n191;
wire n192;
wire n193;
wire n195;
wire n196;
wire n197;
wire n199;
wire n200;
wire n201;
wire n202;
wire n203;
wire n204;
wire n205;
wire n206;
wire n207;
wire n208;
wire n209;
wire n210;
wire n211;
wire n212;
wire n213;
wire n214;
wire n215;
wire n216;
wire n217;
wire n218;
wire n220;
wire n221;
wire n222;
wire n223;
wire n224;
wire n225;
wire n226;
wire n227;
wire n228;
wire n229;
wire n230;
wire n231;
wire n232;
wire n233;
wire n234;
wire n235;
wire n236;
wire n237;
wire n238;
wire n239;
wire n240;
wire n241;
wire n242;
wire n243;
wire n244;
wire n245;
wire n246;
wire n247;
wire n248;
wire n249;
wire n250;
wire n251;
wire n252;
wire n253;
wire n254;
wire n255;
wire n256;
wire n257;
wire n258;
wire n259;
wire n260;
wire n261;
wire n262;
wire n263;
wire n264;
wire n265;
wire n266;
wire n267;
wire n268;
wire n269;
wire n270;
wire n271;
wire n272;
wire n273;
wire n274;
wire n275;
wire n276;
wire n277;
wire n278;
wire n279;
wire n280;
wire n281;
wire n282;
wire n283;
wire n284;
wire n285;
wire n286;
wire n287;
wire n288;
wire n289;
wire n290;
wire n291;
wire n292;
wire n293;
wire n294;
wire n295;
wire n296;
wire n297;
wire n298;
wire n299;
wire n300;
wire n301;
wire n302;
wire n303;
wire n304;
wire n305;
wire n306;
wire n307;
wire n308;
wire n309;
wire n310;
wire n311;
wire n312;
wire n313;
wire n314;
wire n315;
wire n316;
wire n317;
wire n318;
wire n319;
wire n320;
wire n321;
wire n322;
wire n323;
wire n324;
wire n325;
wire n326;
wire n327;
wire n328;
wire n329;
wire n330;
wire n331;
wire n332;
wire n333;
wire n334;
wire n335;
wire n336;
wire n337;
wire n338;
wire n339;
wire n340;
wire n341;
wire n342;
wire n343;
wire n344;
wire n345;
wire n346;
wire n347;
wire n348;
wire n349;
wire n350;
wire n351;
wire n352;
wire n353;
wire n354;
wire n355;
wire n356;
wire n357;
wire n358;
wire n359;
wire n360;
wire n361;
wire n362;
wire n363;
wire n364;
wire n365;
wire n366;
wire n367;
wire n368;
wire n369;
wire n370;
wire n371;
wire n372;
wire n373;
wire n374;
wire n375;
wire n376;
wire n377;
wire n378;
wire n379;
wire n380;
wire n381;
wire n382;
wire n383;
wire n384;
wire n385;
wire n386;
wire n387;
wire n388;
wire n389;
wire n390;
wire n391;
wire n392;
wire n393;
wire n394;
wire n395;
wire n396;
wire n397;
wire n398;
wire n399;
wire n400;
wire n401;
wire n402;
wire n403;
wire n404;
wire n405;
wire n406;
wire n407;
wire n408;
wire n409;
wire n410;
wire n411;
wire n412;
wire n413;
wire n414;
wire n415;
wire n416;
wire n417;
wire n418;
wire n419;
wire n420;
wire n421;
wire n422;
wire n423;
wire n424;
wire n425;
wire n426;
wire n427;
wire n428;
wire n429;
wire n430;
wire n431;
wire n432;
wire n433;
wire n434;
wire n435;
wire n436;
wire n437;
wire n438;
wire n439;
wire n440;
wire n441;
wire n442;
wire n443;
wire n444;
wire n445;
wire n446;
wire n447;
wire n448;
wire n449;
wire n450;
wire n451;
wire n452;
wire n453;
wire n454;
wire n455;
wire n456;
wire n457;
wire n458;
wire n459;
wire n460;
wire n461;
wire n462;
wire n463;
wire n464;
wire n465;
wire n466;
wire n467;
wire n468;
wire n469;
wire n470;
wire n471;
wire n472;
wire n473;
wire n474;
wire n475;
wire n476;
wire n477;
wire n478;
wire n479;
wire n480;
wire n481;
wire n482;
wire n483;
wire n484;
wire n485;
wire n486;
wire n487;
wire n488;
wire n489;
wire n490;
wire n491;
wire n492;
wire n493;
wire n494;
wire n495;
wire n496;
wire n497;
wire n498;
wire n499;
wire n500;
wire n501;
wire n502;
wire n503;
wire n504;
wire n505;
wire n506;
wire n507;
wire n508;
wire n509;
wire n510;
wire n511;
wire n512;
wire n513;
wire n514;
wire n515;
wire n516;
wire n517;
wire n518;
wire n519;
wire n520;
wire n521;
wire n522;
wire n523;
wire n524;
wire n525;
wire n526;
wire n527;
wire n528;
wire n529;
wire n530;
wire n531;
wire n532;
wire n533;
wire n534;
wire n535;
wire n536;
wire n537;
wire n538;
wire n539;
wire n540;
wire n541;
wire n542;
wire n543;
wire n544;
wire n545;
wire n546;
wire n547;
xor (out,n0,n364);
xor (n0,n1,n321);
xor (n1,n2,n166);
xor (n2,n3,n107);
xor (n3,n4,n79);
xor (n4,n5,n45);
or (n5,n6,n37,n44);
and (n6,n7,n18);
and (n7,n8,n11);
and (n8,n9,n10);
xor (n11,n12,n15);
and (n12,n13,n14);
and (n15,n16,n17);
xor (n18,n19,n31);
xor (n19,n20,n21);
and (n20,n12,n15);
xor (n21,n22,n29);
xor (n22,n23,n26);
and (n23,n24,n25);
and (n26,n27,n28);
and (n29,n9,n30);
xor (n31,n32,n35);
xor (n32,n33,n34);
and (n33,n13,n10);
and (n34,n16,n14);
and (n35,n36,n17);
and (n37,n18,n38);
nor (n38,n39,n41);
not (n39,n40);
and (n41,n42,n40);
not (n42,n43);
and (n44,n7,n38);
xor (n45,n46,n65);
xor (n46,n47,n51);
or (n47,n48,n49,n50);
and (n48,n20,n21);
and (n49,n21,n31);
and (n50,n20,n31);
xor (n51,n52,n60);
xor (n52,n53,n57);
or (n53,n54,n55,n56);
and (n54,n23,n26);
and (n55,n26,n29);
and (n56,n23,n29);
nor (n57,n58,n59);
not (n58,n24);
and (n59,n42,n24);
nor (n60,n61,n64);
and (n61,n62,n17);
not (n62,n63);
not (n64,n17);
xor (n65,n66,n76);
xor (n66,n67,n71);
or (n67,n68,n69,n70);
and (n68,n33,n34);
and (n69,n34,n35);
and (n70,n33,n35);
xor (n71,n72,n75);
xor (n72,n73,n74);
and (n73,n13,n30);
and (n74,n16,n10);
and (n75,n36,n14);
xor (n76,n77,n78);
and (n77,n27,n25);
and (n78,n9,n28);
or (n79,n80,n103,n106);
and (n80,n81,n88);
or (n81,n82,n85,n87);
and (n82,n83,n84);
and (n83,n40,n25);
and (n84,n24,n28);
and (n85,n84,n86);
and (n86,n27,n30);
and (n87,n83,n86);
or (n88,n89,n100,n102);
and (n89,n90,n98);
or (n90,n91,n94,n97);
and (n91,n92,n93);
and (n92,n27,n14);
and (n93,n9,n17);
and (n94,n95,n96);
and (n95,n9,n14);
and (n96,n13,n17);
and (n97,n91,n96);
xor (n98,n99,n86);
xor (n99,n83,n84);
and (n100,n98,n101);
xor (n101,n8,n11);
and (n102,n90,n101);
and (n103,n88,n104);
xor (n104,n105,n38);
xor (n105,n7,n18);
and (n106,n81,n104);
or (n107,n108,n136);
and (n108,n109,n111);
xor (n109,n110,n104);
xor (n110,n81,n88);
or (n111,n112,n132,n135);
and (n112,n113,n116);
and (n113,n114,n115);
and (n114,n24,n30);
and (n115,n27,n10);
or (n116,n117,n128,n131);
and (n117,n118,n127);
or (n118,n119,n124,n126);
and (n119,n120,n123);
and (n120,n121,n122);
and (n121,n24,n14);
and (n122,n27,n17);
and (n123,n24,n10);
and (n124,n123,n125);
xor (n125,n92,n93);
and (n126,n120,n125);
xor (n127,n114,n115);
and (n128,n127,n129);
xor (n129,n130,n96);
xor (n130,n91,n95);
and (n131,n118,n129);
and (n132,n116,n133);
xor (n133,n134,n101);
xor (n134,n90,n98);
and (n135,n113,n133);
and (n136,n137,n138);
xor (n137,n109,n111);
or (n138,n139,n161);
and (n139,n140,n142);
xor (n140,n141,n133);
xor (n141,n113,n116);
and (n142,n143,n159);
or (n143,n144,n155,n158);
and (n144,n145,n154);
or (n145,n146,n151,n153);
and (n146,n147,n150);
and (n147,n148,n149);
and (n148,n40,n14);
and (n149,n24,n17);
and (n150,n40,n10);
and (n151,n150,n152);
xor (n152,n121,n122);
and (n153,n147,n152);
and (n154,n40,n30);
and (n155,n154,n156);
xor (n156,n157,n125);
xor (n157,n120,n123);
and (n158,n145,n156);
xor (n159,n160,n129);
xor (n160,n118,n127);
and (n161,n162,n163);
xor (n162,n140,n142);
and (n163,n164,n165);
and (n164,n40,n28);
xor (n165,n143,n159);
xor (n166,n167,n262);
xor (n167,n168,n234);
xor (n168,n169,n201);
or (n169,n170,n195,n200);
and (n170,n171,n179);
and (n171,n172,n174);
and (n172,n173,n10);
xor (n174,n175,n177);
and (n175,n176,n14);
and (n177,n178,n17);
xor (n179,n180,n189);
xor (n180,n181,n182);
and (n181,n175,n177);
xor (n182,n183,n188);
xor (n183,n184,n186);
and (n184,n185,n25);
and (n186,n187,n28);
and (n188,n173,n30);
xor (n189,n190,n193);
xor (n190,n191,n192);
and (n191,n176,n10);
and (n192,n178,n14);
and (n193,n194,n17);
and (n195,n179,n196);
nor (n196,n197,n199);
not (n197,n198);
and (n199,n42,n198);
and (n200,n171,n196);
xor (n201,n202,n220);
xor (n202,n203,n207);
or (n203,n204,n205,n206);
and (n204,n181,n182);
and (n205,n182,n189);
and (n206,n181,n189);
xor (n207,n208,n216);
xor (n208,n209,n213);
or (n209,n210,n211,n212);
and (n210,n184,n186);
and (n211,n186,n188);
and (n212,n184,n188);
nor (n213,n214,n215);
not (n214,n185);
and (n215,n42,n185);
nor (n216,n217,n64);
and (n217,n218,n17);
not (n218,n219);
xor (n220,n221,n231);
xor (n221,n222,n226);
or (n222,n223,n224,n225);
and (n223,n191,n192);
and (n224,n192,n193);
and (n225,n191,n193);
xor (n226,n227,n230);
xor (n227,n228,n229);
and (n228,n176,n30);
and (n229,n178,n10);
and (n230,n194,n14);
xor (n231,n232,n233);
and (n232,n187,n25);
and (n233,n173,n28);
or (n234,n235,n258,n261);
and (n235,n236,n243);
or (n236,n237,n240,n242);
and (n237,n238,n239);
and (n238,n198,n25);
and (n239,n185,n28);
and (n240,n239,n241);
and (n241,n187,n30);
and (n242,n238,n241);
or (n243,n244,n255,n257);
and (n244,n245,n253);
or (n245,n246,n249,n252);
and (n246,n247,n248);
and (n247,n187,n14);
and (n248,n173,n17);
and (n249,n250,n251);
and (n250,n173,n14);
and (n251,n176,n17);
and (n252,n246,n251);
xor (n253,n254,n241);
xor (n254,n238,n239);
and (n255,n253,n256);
xor (n256,n172,n174);
and (n257,n245,n256);
and (n258,n243,n259);
xor (n259,n260,n196);
xor (n260,n171,n179);
and (n261,n236,n259);
or (n262,n263,n291);
and (n263,n264,n266);
xor (n264,n265,n259);
xor (n265,n236,n243);
or (n266,n267,n287,n290);
and (n267,n268,n271);
and (n268,n269,n270);
and (n269,n185,n30);
and (n270,n187,n10);
or (n271,n272,n283,n286);
and (n272,n273,n282);
or (n273,n274,n279,n281);
and (n274,n275,n278);
and (n275,n276,n277);
and (n276,n185,n14);
and (n277,n187,n17);
and (n278,n185,n10);
and (n279,n278,n280);
xor (n280,n247,n248);
and (n281,n275,n280);
xor (n282,n269,n270);
and (n283,n282,n284);
xor (n284,n285,n251);
xor (n285,n246,n250);
and (n286,n273,n284);
and (n287,n271,n288);
xor (n288,n289,n256);
xor (n289,n245,n253);
and (n290,n268,n288);
and (n291,n292,n293);
xor (n292,n264,n266);
or (n293,n294,n316);
and (n294,n295,n297);
xor (n295,n296,n288);
xor (n296,n268,n271);
and (n297,n298,n314);
or (n298,n299,n310,n313);
and (n299,n300,n309);
or (n300,n301,n306,n308);
and (n301,n302,n305);
and (n302,n303,n304);
and (n303,n198,n14);
and (n304,n185,n17);
and (n305,n198,n10);
and (n306,n305,n307);
xor (n307,n276,n277);
and (n308,n302,n307);
and (n309,n198,n30);
and (n310,n309,n311);
xor (n311,n312,n280);
xor (n312,n275,n278);
and (n313,n300,n311);
xor (n314,n315,n284);
xor (n315,n273,n282);
and (n316,n317,n318);
xor (n317,n295,n297);
and (n318,n319,n320);
and (n319,n198,n28);
xor (n320,n298,n314);
or (n321,n322,n325,n363);
and (n322,n323,n324);
xor (n323,n137,n138);
xor (n324,n292,n293);
and (n325,n324,n326);
or (n326,n327,n330,n362);
and (n327,n328,n329);
xor (n328,n162,n163);
xor (n329,n317,n318);
and (n330,n329,n331);
or (n331,n332,n335,n361);
and (n332,n333,n334);
xor (n333,n164,n165);
xor (n334,n319,n320);
and (n335,n334,n336);
or (n336,n337,n342,n360);
and (n337,n338,n340);
xor (n338,n339,n156);
xor (n339,n145,n154);
xor (n340,n341,n311);
xor (n341,n300,n309);
and (n342,n340,n343);
or (n343,n344,n349,n359);
and (n344,n345,n347);
xor (n345,n346,n152);
xor (n346,n147,n150);
xor (n347,n348,n307);
xor (n348,n302,n305);
and (n349,n347,n350);
or (n350,n351,n354,n358);
and (n351,n352,n353);
xor (n352,n148,n149);
xor (n353,n303,n304);
and (n354,n353,n355);
and (n355,n356,n357);
and (n356,n40,n17);
and (n357,n198,n17);
and (n358,n352,n355);
and (n359,n345,n350);
and (n360,n338,n343);
and (n361,n333,n336);
and (n362,n328,n331);
and (n363,n323,n326);
xor (n364,n365,n489);
xor (n365,n366,n461);
xor (n366,n367,n428);
xor (n367,n368,n377);
and (n368,n369,n373);
nor (n369,n370,n372);
not (n370,n371);
xor (n371,n40,n198);
and (n372,n42,n371);
and (n373,n374,n25);
xor (n374,n375,n376);
xor (n375,n24,n185);
and (n376,n40,n198);
or (n377,n378,n425,n427);
and (n378,n379,n406);
and (n379,n380,n391);
and (n380,n381,n10);
xor (n381,n382,n383);
xor (n382,n9,n173);
or (n383,n384,n385,n390);
and (n384,n27,n187);
and (n385,n187,n386);
or (n386,n387,n388,n389);
and (n387,n24,n185);
and (n388,n185,n376);
and (n389,n24,n376);
and (n390,n27,n386);
xor (n391,n392,n399);
and (n392,n393,n14);
xor (n393,n394,n395);
xor (n394,n13,n176);
or (n395,n396,n397,n398);
and (n396,n9,n173);
and (n397,n173,n383);
and (n398,n9,n383);
and (n399,n400,n17);
xor (n400,n401,n402);
xor (n401,n16,n178);
or (n402,n403,n404,n405);
and (n403,n13,n176);
and (n404,n176,n395);
and (n405,n13,n395);
xor (n406,n407,n416);
xor (n407,n408,n409);
and (n408,n392,n399);
xor (n409,n410,n415);
xor (n410,n411,n414);
and (n411,n412,n28);
xor (n412,n413,n386);
xor (n413,n27,n187);
and (n414,n381,n30);
and (n415,n393,n10);
xor (n416,n417,n418);
and (n417,n400,n14);
and (n418,n419,n17);
xor (n419,n420,n421);
xor (n420,n36,n194);
or (n421,n422,n423,n424);
and (n422,n16,n178);
and (n423,n178,n402);
and (n424,n16,n402);
and (n425,n406,n426);
xor (n426,n369,n373);
and (n427,n379,n426);
xor (n428,n429,n440);
xor (n429,n430,n434);
or (n430,n431,n432,n433);
and (n431,n408,n409);
and (n432,n409,n416);
and (n433,n408,n416);
xor (n434,n435,n439);
or (n435,n436,n437,n438);
and (n436,n411,n414);
and (n437,n414,n415);
and (n438,n411,n415);
and (n439,n417,n418);
xor (n440,n441,n456);
xor (n441,n442,n445);
nor (n442,n443,n444);
not (n443,n374);
and (n444,n42,n374);
xor (n445,n446,n449);
xor (n446,n447,n448);
and (n447,n400,n10);
and (n448,n419,n14);
and (n449,n450,n17);
xor (n450,n451,n452);
xor (n451,n63,n219);
or (n452,n453,n454,n455);
and (n453,n36,n194);
and (n454,n194,n421);
and (n455,n36,n421);
xor (n456,n457,n460);
xor (n457,n458,n459);
and (n458,n412,n25);
and (n459,n381,n28);
and (n460,n393,n30);
or (n461,n462,n485,n488);
and (n462,n463,n470);
or (n463,n464,n467,n469);
and (n464,n465,n466);
and (n465,n371,n25);
and (n466,n374,n28);
and (n467,n466,n468);
and (n468,n412,n30);
and (n469,n465,n468);
or (n470,n471,n482,n484);
and (n471,n472,n480);
or (n472,n473,n476,n479);
and (n473,n474,n475);
and (n474,n412,n14);
and (n475,n381,n17);
and (n476,n477,n478);
and (n477,n381,n14);
and (n478,n393,n17);
and (n479,n473,n478);
xor (n480,n481,n468);
xor (n481,n465,n466);
and (n482,n480,n483);
xor (n483,n380,n391);
and (n484,n472,n483);
and (n485,n470,n486);
xor (n486,n487,n426);
xor (n487,n379,n406);
and (n488,n463,n486);
or (n489,n490,n518);
and (n490,n491,n493);
xor (n491,n492,n486);
xor (n492,n463,n470);
or (n493,n494,n514,n517);
and (n494,n495,n498);
and (n495,n496,n497);
and (n496,n374,n30);
and (n497,n412,n10);
or (n498,n499,n510,n513);
and (n499,n500,n509);
or (n500,n501,n506,n508);
and (n501,n502,n505);
and (n502,n503,n504);
and (n503,n374,n14);
and (n504,n412,n17);
and (n505,n374,n10);
and (n506,n505,n507);
xor (n507,n474,n475);
and (n508,n502,n507);
xor (n509,n496,n497);
and (n510,n509,n511);
xor (n511,n512,n478);
xor (n512,n473,n477);
and (n513,n500,n511);
and (n514,n498,n515);
xor (n515,n516,n483);
xor (n516,n472,n480);
and (n517,n495,n515);
and (n518,n519,n520);
xor (n519,n491,n493);
or (n520,n521,n543);
and (n521,n522,n524);
xor (n522,n523,n515);
xor (n523,n495,n498);
and (n524,n525,n541);
or (n525,n526,n537,n540);
and (n526,n527,n536);
or (n527,n528,n533,n535);
and (n528,n529,n532);
and (n529,n530,n531);
and (n530,n371,n14);
and (n531,n374,n17);
and (n532,n371,n10);
and (n533,n532,n534);
xor (n534,n503,n504);
and (n535,n529,n534);
and (n536,n371,n30);
and (n537,n536,n538);
xor (n538,n539,n507);
xor (n539,n502,n505);
and (n540,n527,n538);
xor (n541,n542,n511);
xor (n542,n500,n509);
and (n543,n544,n545);
xor (n544,n522,n524);
and (n545,n546,n547);
and (n546,n371,n28);
xor (n547,n525,n541);
endmodule
